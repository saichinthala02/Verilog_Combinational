module mux161(i,s,y);
  input [15:0]i;
  input [3:0]s;
  output reg y;

  always@(s)begin
    case(s)
      4'b0000 : y=i[0];
      4'b0001 : y=i[1];
      4'b0010 : y=i[2];
      4'b0011 : y=i[3];
      4'b0100 : y=i[4];
      4'b0101 : y=i[5];
      4'b0110 : y=i[6];
      4'b0111 : y=i[7];
      4'b1000 : y=i[8];
      4'b1001 : y=i[9];
      4'b1010 : y=i[10];
      4'b1011 : y=i[11];
      4'b1100 : y=i[12];
      4'b1101 : y=i[13];
      4'b1110 : y=i[14];
      4'b1111 : y=i[15];
      default : y=4'bxxxx;
    endcase
  end
endmodule 

module top;
  reg [15:0]i;
  reg [3:0]s;
  wire y;
  mux161 dut(i,s,y);
  initial begin
    $display("------------------------------------");
    $display("------------> 16x1 MUX <------------");
    $display("------------------------------------");
    $display("|        i         |   s  |  Yout |");
    $display("------------------------------------");
    repeat(10)begin
      {i,s}=$random;
      #2 $display("| %b | %b |   %b   |",i,s,y);
    end
    $display("------------------------------------");
  end
endmodule
/* Output:-
# Start time: 11:21:39 on Oct 04,2025
# Loading work.top
# Loading work.mux161
# ------------------------------------
# ------------> 16x1 MUX <------------
# ------------------------------------
# |        i         |   s  |  Yout |
# ------------------------------------
# | 0101001101010010 | 0100 |   1   |
# | 1001010111101000 | 0001 |   0   |
# | 0100110101100000 | 1001 |   0   |
# | 0000010101100110 | 0011 |   0   |
# | 1001011110110000 | 1101 |   0   |
# | 1111100110011000 | 1101 |   0   |
# | 0010100001000110 | 0101 |   0   |
# | 0111010100100001 | 0010 |   0   |
# | 0011111000110000 | 0001 |   0   |
# | 0111110011010000 | 1101 |   1   |
# ------------------------------------
*/
